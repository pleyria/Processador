module Bin2BCD (clock, bin, start, bcd);

input clock, start;
input [15:0] bin;

output [19:0] bcd;

// aliases para os estados
parameter s_INATIVO = 3'b000;
parameter s_SHIFT = 3'b001;
parameter s_VERIFICA_SHIFT = 3'b010;
parameter s_SOMA = 3'b011;
parameter s_VERIFICA_DIGITO_DECIMAL = 3'b100;
parameter s_FIM = 3'b101;

// registrador para o estado da maquina de estados
reg [2:0] estado;

// registrador para a saida em BCD
reg [19:0] r_bcd;

// registrador para a entrada em binario
reg [15:0] r_bin;

// registrador para o digito decimal
reg [4:0] digito_decimal;

// registrador para iteracoes
reg [3:0] i;

// conexao para o digito atual bcd analisado
wire [3:0] digito_BCD;

assign digito_BCD = r_bcd[(digito_decimal*4) +: 4];
assign bcd = r_bcd;

initial begin
	estado = s_INATIVO;
	i = 0;
	digito_decimal = 0;
end

always @ (posedge clock) begin

	case (estado)

		// fica no estado inicial ate receber o sinal de start
		s_INATIVO: begin
			if (start) begin
				r_bin <= bin;
				estado <= s_SHIFT;
				r_bcd <= 0;
			end
			else begin
				estado <= s_INATIVO;
			end
		end

		// Faz o shift para bcd ate o ultimo bit binario
		s_SHIFT: begin
			r_bcd <= r_bcd << 1;
			r_bcd[0] <= r_bin[15];
			r_bin <= r_bin << 1;
			estado <= s_VERIFICA_SHIFT;
		end

		// Verifica se acabou o shift do binario
		s_VERIFICA_SHIFT: begin
			if (i == 4'd15) begin
				i <= 0;
				estado <= s_FIM;
			end
			else begin
				i <= i + 4'b1;
				estado <= s_SOMA;
			end
		end

		// Verifica se precisa somar 3 no bcd
		s_SOMA: begin
			if (digito_BCD > 4) begin
				r_bcd[(digito_decimal*4) +: 4] <= digito_BCD + 20'd3;
			end
			estado <= s_VERIFICA_DIGITO_DECIMAL;
		end

		// Verifica se somou 3 a todos os digitos
		s_VERIFICA_DIGITO_DECIMAL: begin
			if (digito_decimal == 5'd4) begin
				digito_decimal <= 0;
				estado <= s_SHIFT;
			end
			else begin
				digito_decimal <= digito_decimal + 5'b1;
				estado <= s_SOMA;
			end
		end

		// Fim da decodificacao
		s_FIM:
			estado <= s_INATIVO;

		default:
			estado <= s_INATIVO;

	endcase
	
end

endmodule
